----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Xandão e Xandona
-- 
-- Create Date:    14:38:16 11/25/2025 
-- Design Name: 
-- Module Name:    xandinho - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity xandinho is
port(
	clk, inicializar : in std_logic;
	debugEndereco : in std_logic_vector (9 downto 2);
	debugPalavra : out std_logic_vector (9 downto 2)
);
end xandinho;

architecture Behavioral of xandinho is
--pc
	component pc is
		port(
			ini, clk : in std_logic;
			entrada : in std_logic_vector(31 downto 0);
			saida : out std_logic_vector(31 downto 0)
		);
		end component;
--memInstrucoes
	component memInstrucoes is
	port (
		Endereco : in std_logic_vector(31 downto 0);
		Palavra : out std_logic_vector(31 downto 0)
	);
end component;
	
--unidade_controle
	component unidade_controle is
    port(
        op_uc : in std_logic_vector(5 downto 0); 
        ALU_op_uc : out std_logic_vector (1 downto 0); 
        reg_write, reg_dst, ALU_src, branch, mem_write, mem_toReg, jump, mem_read : out std_logic
    );
end component;
--mux2
	component mux2 is
	port(
		A, B, s: in std_logic;
		resultado : out std_logic
	);
end component;
--banco_registradores
	component banco_registradores is
    port(
        clk, escreverReg : in std_logic;
        dadoEscrita : in std_logic_vector (31 downto 0); -- alexandre - mudei pra down to 
        endEscrita : in std_logic_vector (4 downto 0); -- mudei

        endL1 : in std_logic_vector(4 downto 0);
        endL2 : in std_logic_vector(4 downto 0);

        dadoL1 : out std_logic_vector(31 downto 0); 
        dadoL2 : out std_logic_vector(31 downto 0)
    );
end component;

--extensor_sinal
	component extensor_sinal is
    port(
        entrada_16 : in std_logic_vector (15 downto 0);
        saida_32   : out std_logic_vector (31 downto 0)
    );
end component;
--uc_ula
	component uc_ula is
    port(
    ALU_op : in std_logic_vector (1 downto 0);
    funct : in std_logic_vector (5 downto 0);
    Ainverte, Binverte : out std_logic;
    operacao : out std_logic_vector (1 downto 0)
    );
end component;
--ula_32
	component ula_32 is
	port(
		a : in std_logic_vector (31 downto 0); -- mudei pra downto
        b : in std_logic_vector (31 downto 0); -- mudei pra downto
		Ainverte, Binverte : in std_logic;
		op : in std_logic_vector(1 downto 0);--alexandre - corrigi auqi pra um vetor de 2 
		result : out std_logic_vector (31 downto 0); -- mudei pra downto
		zero : out std_logic
	);
end component;
--memDados
	component memDados is
	port (
		DadoLido : out std_logic_vector (31 downto 0);
		DadoEscrita : in std_logic_vector (31 downto 0);
		Endereco : in std_logic_vector (31 downto 0);
		EscreverMem : in std_logic;
		Clock : in std_logic;
		LerMem : in std_logic;
		DebugEndereco : in std_logic_vector(31 downto 0);
		DebugPalavra : out std_logic_vector(31 downto 0));
end component;
--somador
	component somador is
	port(
	A, B : in std_logic;
	vai1, saida : out std_logic
	);
end component;
--somador completo
	component somador_completo is
	port(
	A, B, vem1 : in std_logic;
	vai1, resultado : out std_logic
	);
end component;
--deslocador_2
	component deslocador_2 is
    port(
        entrada_32 : in std_logic_vector (31 downto 0);
        saida_32   : out std_logic_vector (31 downto 0)
    );
end component;
	--signal 1 :
	signal saidaPC : std_logic_vector(31 downto 0);
	--signal 2 :
	signal saidaMemoInstru : std_logic_vector(31 downto 0);
	--signal 3 :
	signal saidaUC_regDst : std_logic;
	--signal 4:
	signal saidaMuxA_bancoReg : std_logic_vector(4 downto 0);
	--signal 5:
	signal saidaMuxC_writeData_bancoReg : std_logic_vector(31 downto 0);
	--signal 6:
	signal saidaUC_regWrite : std_logic;
	--signal 7:
	signal saidaData1_ULA : std_logic_vector(31 downto 0);
	--signal 8:
	signal saidaData2 : std_logic_vector(31 downto 0);
	--signal 9:
	signal saidaExtSinal_deslocA : std_logic_vector(31 downto 0);
	--signal 10:
	signal saidaUC_muxB : std_logic;
	--signal 11:
	signal saidaMuxB_ULA : std_logic_vector(31 downto 0);
	--signal 12:
	signal saidaUC_UCula : std_logic;
	--signal 13:
	signal saidaUCula_ULA : std_logic_vector(1 downto 0);-- mais de 1 sinal
	--signal 14:
	signal saidaZeroULA_and : std_logic;
	--signal 15:
	signal saidaULA : std_logic_vector(31 downto 0);
	--signal 16:
	signal saidaUC_memWrite : std_logic;
	--signal 17:
	signal saidaDataMem_muxC : std_logic_vector(31 downto 0);
	--signal 18:
	signal saidaUC_memRead : std_logic;
	--signal 19:
	signal saidaUC_memtoReg : std_logic;
	--signal 20: (esse n tem)
	--signal
	--signal 21:
	signal saidaSomadorA : std_logic_vector(31 downto 0);--acho q esse aqui vai ter q ser vetor
	--signal 22:
	signal saidaDeslocB_muxE : std_logic_vector(31 downto 0);--atecnao pra esse aqui, ele meio q se junta com esse de cima
	--signal 23:
	signal saidaDeslocA_somadorB : std_logic_vector(31 downto 0);
	--signal 24:
	signal saidaSomadorB_muxD : std_logic_vector(31 downto 0);
	--signal 25:
	signal saidaUC_branch : std_logic;
	--signal 26:
	signal saidaAnd_muxD : std_logic;
	--signal 27:
	signal saidaMuxD_muxE : std_logic_vector(31 downto 0);
	--signal 28:
	signal saidaUC_jump : std_logic;
	--signal 29:
	signal saidaMuxE_pc : std_logic_vector(31 downto 0);

	
begin
	--port map do pc:
	PC_reg: pc port map(
		ini => inicializar,
		clk => clk,
		entrada => saidaMuxE_pc, -- 29
		saida => saidaPC -- 1
		);

	-- port map memoria de instrucao
	memoria_inst: memInstrucoes port map(
		Endereco => saidaPC,
		Palavra => saidaMemoInstru -- fio 2
    	);

	-- port map unidade de controle
	uc_principal: unidade_controle port map(
		op_uc => saidaMemoInstru(31 downto 26), 
	    ALU_op_uc => ALU_op_control,
	    reg_write => saidaUC_regWrite,
	    reg_dst => saidaUC_regDst,
	    ALU_src => saidaUC_muxB,
	    branch => saidaUC_branch,
	    mem_write => saidaUC_memWrite,
	    mem_toReg => saidaUC_memtoReg,
	    jump => saidaUC_jump,
	    mem_read => saidaUC_memRead
		);

	--port map muxA
	mux_A : mux2 port map(
		A => saidaMemoInstru(20 downto 16),
		B => saidaMemoInstru(15 downto 11),
		s => saidaUC_regDst, -- fio 3
		resultado => saidaMuxA_bancoReg
		);

	-- port map unidade de controla da ula
	UC_ula : uc_ula port map(
		ALU_op => saidaUC_UCula, --fio 12
		operacao => saidaUCula_ULA, -- fio 13, obs: na imagemd e caminho da dados fala "mais de 1 sinal"
		funct => saidaMemoInstru(5 downto 0)
		--Ainverte ?
		--Binverte ?
		);

	--port map extensor de sinal
	extensor_de_sinal is extensor_sinal port map(
		entrada_16 => saidaMemoInstru(15 downto 0),
		saida_32 => saidaExtSinal_deslocA -- fio 9
		);
	

	--port map banco de registradores
	banco_de_resgistradores : banco_registradores port map(
		clk => clk;
		endL1 => saidaMemoInstru(25 downto 21),
		endL2 => saidaMemoInstru(25 downto 21),
		escreverReg => saidaMuxA_bancoReg, --fio 4
		dadoEscrita => saidaMuxC_writeData_bancoReg -- fio5
		dadoL1 => saidaData1_ULA -- fio 7
		dadoL2 => 	saidaData2 -- aqui tem q ver pq ele vai pra dois lugares
	    );

	--port map muxB
	mux_B : mux2 port map(
		A => saidaData1_ULA, -- fio 8
		B => saidaExtSinal_deslocA, -- fio 9, tem q ver aqui pq esse fio vai pra 2 lugares
		s => saidaUC_muxB, --fio 10
		resultado => saidaMuxB_ULA -- fio 11
		);

	--port map ula
	ula_principal : ula_32 port map(
		a => saidaData1_ULA,  -- fio 7
		b => saidaMuxB_ULA, -- fio 11
		op = > saidaUCula_ULA, -- fio 13
		zero => saidaZeroULA_and, -- fio 14
		result => saidaULA, -- fio 15, tem q ver aqui pq ele vai pra dois lugares diferentes
		--Ainverte e Binverte??
		);

	-- port map memoria de dados
	memoria_de_dados : memDados port map(
		DadoLido => saidaULA, -- fio 15, tem q ver aqui pq esse fio vai pra 2 lugares7
		DadoEscrita => saidaData2, -- fio 8,  tem q ver aqui pq esse fio vai pra 2 lugares7
		Clock => clk,
		LerMem => saidaDataMem_muxC, -- fio 17
		--OS FIOS 16 E 18 VAO PRA ALGUM LUGAR AQUI
		Endereco => 
		EscreverMem =>
		DebugEndereco =>
		DebugPalavra =>
		);

	--port map mux c
	mux_C : mux2 port map(
		B => saidaDataMem_muxC, -- fio 17
		A => saidaULA, -- fio 15, tem q ver aqui pq esse fio vai pra 2 lugares
		s => saidaUC_memtoReg, -- fio 19
		resultado => saidaMuxC_writeData_bancoReg -- fio 5
	    );

	--port map somador A
	somador_A is somador port map(
		
	
		);

	-- port map deslocador B
	deslocador_B is delocador_2 port map(
		entrada_32 => saidaMemoInstru(25 downto 0),
		saida_32 => saidaDeslocB_muxE -- fio 22
		);

	-- port map deslocador A 
	deslocador_B is delocador_2 port map(
		entrada_32 => saidaExtSinal_deslocA,
		saida_32 => saidaDeslocA_somadorB -- fio 23
		);

	--port map muxD
	mux_D : mux2 port map(
		A => saidaSomadorA, -- FIO 21
		B => saidaSomadorB_muxD, -- FIO 24
		s=> saidaAnd_muxD, -- fio 26
		resultado => saidaMuxD_muxE -- fio 27
		);

	--port map muxE
	mux_E : mux2 port map(
		B => saidaDeslocB_muxE, -- FIO 22, SE ATENTAR AQUI PQ TEM QUE FAZER SLICE NESSE FIO
		A => saidaMuxD_muxE, -- FIO 27
		s=> saidaUC_jump, -- fio 28
		resultado => saidaMuxE_pc -- fio 29
		);

	
end Behavioral;

